library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
	type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType : TPicoType := pbt3 ;
	function ADDRSIZE return natural ;
	function INSTSIZE return natural ;
	function JADDRSIZE return natural ;
	function JDATASIZE return natural ;
end package ;

package body constants is
	function ADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 10 ;
		when pbt3 => return 10 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function INSTSIZE return natural is 
	begin
		case PicoType is
		when pbtI => return 16 ;
		when pbtII => return 18 ;
		when pbt3 => return 18 ;
		when pbtS => return 18 ;
		end case ;
	end ;
	function JADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 9 ;
		when pbtII => return 11 ;
		when pbt3 => return 11 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function JDATASIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 9 ;
		when pbt3 => return 9 ;
		when pbtS => return 20 ;
		end case ;
	end ;
end package body ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;

use work.constants.all;

entity memoria is
    port ( 
        clk : in std_logic ;
        reset : out std_logic ;
        address : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity memoria ;

architecture mix of memoria is
    component jtag_shifter is
        port ( 
			clk : in std_logic ;
			user1 : out std_logic ;
            write : out std_logic ;
            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
        ) ;
    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18 : if (PicoType = pbtII) or (PicoType = pbt3) generate
	    attribute INIT_00 of bram : label is "0000000000000000000000008001C401E4FF50082401440040021BB0C001F440" ;
	    attribute INIT_01 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_02 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_07 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_08 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_09 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_0F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_10 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_11 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_12 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_13 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_14 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_15 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_16 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_17 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_18 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_19 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_35 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "4004000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_00 of bram : label is "00000000000000000000000000000000000000000000000000000000000E34CC" ;
	    attribute INITP_01 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_02 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "C000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"0000000000000000000000008001C401E4FF50082401440040021BB0C001F440",
	            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"4004000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"00000000000000000000000000000000000000000000000000000000000E34CC",
	            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )
	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk,
	            ADDRB => address,

DOB => instruction( 18 - 3 downto 0 ),-- OJO INSTSIZE =18
DOPB => instruction( 18 - 1 downto 18 - 2 ),-- INSTSIZE = 18
DIA => jdata( 9 - 2 downto 0 ),	 -- OJO JDATASIZE = 9
DIPA => jdata( 9 - 1 downto 9 - 1 ), -- OJO JDATASIZE = 9

	            --DOB => instruction( INSTSIZE - 3 downto 0 ),
	            --DOPB => instruction( INSTSIZE - 1 downto INSTSIZE - 2 ),
	            --DIA => jdata( JDATASIZE - 2 downto 0 ),
	            --DIPA => jdata( JDATASIZE - 1 downto JDATASIZE - 1 ),
	            
					ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	I16 : if PicoType = pbtI generate
		attribute INIT_00 of bram : label is "0000000000000000000000008001C401E4FF50082401440040021BB0C001F440" ;
		attribute INIT_01 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_02 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB4_S8_S16
	        generic map (
	            INIT_00 => X"0000000000000000000000008001C401E4FF50082401440040021BB0C001F440",
	            INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIB => "0000000000000000",  
				ENB => '1', 
				WEB => '0',
				RSTB =>	'0',
				CLKB => clk,
				ADDRB => address,
				DOB => instruction( INSTSIZE - 1 downto 0 ),  
				DIA => jdata( JDATASIZE - 1 downto 0 ),   
				ENA => juser1, 
				WEA => jwrite,
				RSTA => '0',
				CLKA => clk,
				ADDRA => jaddr,
				DOA => open  
			) ; 
	end generate ;

	I20 : if PicoType = pbtS generate
		attribute INIT_00 of ram_1 : label is "0000000000000000000000000000000000000000000000000000003203103030" ;
		attribute INIT_01 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_02 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_03 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_04 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_05 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_1 : label is "3000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_2 : label is "0000000000000000000000000000000000000000000000000000008CE52441CF" ;
		attribute INIT_01 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_02 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_03 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_04 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_05 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_2 : label is "4000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000440440B04" ;
		attribute INIT_01 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_02 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_03 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_04 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_05 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_4 : label is "00000000000000000000000000000000000000000000000000000000F0000B04" ;
		attribute INIT_01 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_02 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_03 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_04 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_05 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_5 : label is "00000000000000000000000000000000000000000000000000000011F8102010" ;
		attribute INIT_01 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_02 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_03 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_04 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_05 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_5 : label is "4000000000000000000000000000000000000000000000000000000000000000" ;

		signal data_out : std_logic_vector( 3 downto 0 ) ;
	begin
	    ram_1 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000003203103030",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"3000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => data_out,  
DIB => jdata( 11 downto 9 - 1 ), -- OJO JDATASIZE = 9 Y LOS DI VUELTA  ademas cambiamos el tama�o a 4 bits

				--DIB => jdata( JDATASIZE - 1 downto 16 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
			-- loose top 2 bits
			instruction( 17 downto 16 ) <= data_out( 1 downto 0 ) ;

	    ram_2 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000008CE52441CF",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"4000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 15 downto 12 ),  
				DIB => jdata( 15 downto 12 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_3 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000440440B04",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 11 downto 8 ),  
				DIB => jdata( 11 downto 8 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_4 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"00000000000000000000000000000000000000000000000000000000F0000B04",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 7 downto 4 ),  
				DIB => jdata( 7 downto 4 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_5 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"00000000000000000000000000000000000000000000000000000011F8102010",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"4000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 3 downto 0 ),  
				DIB => jdata( 3 downto 0 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
	end generate ;

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture mix ;
