--------------------------------------------------------------------------------
-- Company: DSI / FCEIA / UNR 
-- Engineer: Curso s�ntesis de sistemas digitales en FPGA - 2016
--
-- Create Date:    10:16:12 05/10/16
-- Design Name:    
-- Module Name:    compara - Behavioral
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description: comparador de n�meros de 4 bits
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments: Modificar para que trabaje con n�meros positivos sin signo.
-- 
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity compara is
    Port ( a : in std_logic_vector(3 downto 0);
           b : in std_logic_vector(3 downto 0);
           mayor: out std_logic);  
end compara;

architecture Behavioral of compara is

begin
mayor <= '1' when a > b else '0';
end Behavioral;
