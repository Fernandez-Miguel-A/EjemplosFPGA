library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
	type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType : TPicoType := pbt3 ;
	function ADDRSIZE return natural ;
	function INSTSIZE return natural ;
	function JADDRSIZE return natural ;
	function JDATASIZE return natural ;
end package ;

package body constants is
	function ADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 10 ;
		when pbt3 => return 10 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function INSTSIZE return natural is 
	begin
		case PicoType is
		when pbtI => return 16 ;
		when pbtII => return 18 ;
		when pbt3 => return 18 ;
		when pbtS => return 18 ;
		end case ;
	end ;
	function JADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 9 ;
		when pbtII => return 11 ;
		when pbt3 => return 11 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function JDATASIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 9 ;
		when pbt3 => return 9 ;
		when pbtS => return 20 ;
		end case ;
	end ;
end package body ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;

use work.constants.all;

entity memoria is
    port ( 
        clk : in std_logic ;
        reset : out std_logic ;
        address : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity memoria ;

architecture mix of memoria is
    component jtag_shifter is
        port ( 
			clk : in std_logic ;
			user1 : out std_logic ;
            write : out std_logic ;
            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
        ) ;
    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18 : if (PicoType = pbtII) or (PicoType = pbt3) generate
	    attribute INIT_00 of bram : label is "C00000BF00BFC00154174900501749FFC000FAA009FFF7700F20001A00EEC000" ;
	    attribute INIT_01 of bram : label is "00BF00DD50234500450406004007CA01C0010AFF4017EAFF54174900501649FF" ;
	    attribute INIT_02 of bram : label is "860100CE051800BA00BA00BA060100BF00BF00BF00BF00BF00BF401B860100BF" ;
	    attribute INIT_03 of bram : label is "00DD052000DD052000DD052000DD05200104051000BF00BF00BF00BF542A4610" ;
	    attribute INIT_04 of bram : label is "00DD052000DD052000DD053A00DD057300DD056F00DD057400DD056100DD0544" ;
	    attribute INIT_05 of bram : label is "A00000DD0520A00054534610860100CE051C00BA00BA00BA00BA060100DD0520" ;
	    attribute INIT_06 of bram : label is "47615874475B587347415874473A58734730157001048F010F2E5864452F15F0" ;
	    attribute INIT_07 of bram : label is "408109FF5C80480AA80F187054804830A8F018700AFF00DD053F5874477B5873" ;
	    attribute INIT_08 of bram : label is "090F0098408F00DD053F01048F010F2E5889452F15F0588E4C0A1C7080000900" ;
	    attribute INIT_09 of bram : label is "C53040A500A6589F450A15C0010415F040811A709780070608075894270FF880" ;
	    attribute INIT_0A of bram : label is "A00054ADC001000BA0000F20001A0104051000EEA0000F2F58A54F2F8F0100DD" ;
	    attribute INIT_0B of bram : label is "037DA00054BBC30100B50314A00054B6C20100B00219A00054B1C10100AC0128" ;
	    attribute INIT_0C of bram : label is "A4F01450A00000C4C440A4F8A000C440E40100ACC440E401A00054C0C30100B5" ;
	    attribute INIT_0D of bram : label is "C40CA4F01450A000C44004F000B000CA0406040604060407145000AC00CAC408" ;
	    attribute INIT_0E of bram : label is "043000BAA000C44004F000B000C4C4400406040604070407145000AC00C4C440" ;
	    attribute INIT_0F of bram : label is "050100CE050C00CE050600CE052800B000CA042000B000CA00B500CA00BA00CA" ;
	    attribute INIT_10 of bram : label is "18704701A00000CEC5C0A50FA00000CEC580A50F510A2510A00000B500B500CE" ;
	    attribute INIT_11 of bram : label is "00000000000000000000000000000000000000000000000040605082A880A77F" ;
	    attribute INIT_12 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_13 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_14 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_15 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_16 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_17 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_18 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_19 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_35 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "410E000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_00 of bram : label is "CD0D033777774D34B2D73FCCCCCCCCCCCCCCCFFD73F3FFF7FD0ECCDDFFDDC03F" ;
	    attribute INITP_01 of bram : label is "3333CFFF3A3EAA3E028FAA3C0B8A38B72DCB72DCB48F38D73F4CC6B43F34D34C" ;
	    attribute INITP_02 of bram : label is "000000000000000000000000000000000000000000000000000000F00B0B0DBF" ;
	    attribute INITP_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "C000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"C00000BF00BFC00154174900501749FFC000FAA009FFF7700F20001A00EEC000",
	            INIT_01 => X"00BF00DD50234500450406004007CA01C0010AFF4017EAFF54174900501649FF",
	            INIT_02 => X"860100CE051800BA00BA00BA060100BF00BF00BF00BF00BF00BF401B860100BF",
	            INIT_03 => X"00DD052000DD052000DD052000DD05200104051000BF00BF00BF00BF542A4610",
	            INIT_04 => X"00DD052000DD052000DD053A00DD057300DD056F00DD057400DD056100DD0544",
	            INIT_05 => X"A00000DD0520A00054534610860100CE051C00BA00BA00BA00BA060100DD0520",
	            INIT_06 => X"47615874475B587347415874473A58734730157001048F010F2E5864452F15F0",
	            INIT_07 => X"408109FF5C80480AA80F187054804830A8F018700AFF00DD053F5874477B5873",
	            INIT_08 => X"090F0098408F00DD053F01048F010F2E5889452F15F0588E4C0A1C7080000900",
	            INIT_09 => X"C53040A500A6589F450A15C0010415F040811A709780070608075894270FF880",
	            INIT_0A => X"A00054ADC001000BA0000F20001A0104051000EEA0000F2F58A54F2F8F0100DD",
	            INIT_0B => X"037DA00054BBC30100B50314A00054B6C20100B00219A00054B1C10100AC0128",
	            INIT_0C => X"A4F01450A00000C4C440A4F8A000C440E40100ACC440E401A00054C0C30100B5",
	            INIT_0D => X"C40CA4F01450A000C44004F000B000CA0406040604060407145000AC00CAC408",
	            INIT_0E => X"043000BAA000C44004F000B000C4C4400406040604070407145000AC00C4C440",
	            INIT_0F => X"050100CE050C00CE050600CE052800B000CA042000B000CA00B500CA00BA00CA",
	            INIT_10 => X"18704701A00000CEC5C0A50FA00000CEC580A50F510A2510A00000B500B500CE",
	            INIT_11 => X"00000000000000000000000000000000000000000000000040605082A880A77F",
	            INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"410E000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"CD0D033777774D34B2D73FCCCCCCCCCCCCCCCFFD73F3FFF7FD0ECCDDFFDDC03F",
	            INITP_01 => X"3333CFFF3A3EAA3E028FAA3C0B8A38B72DCB72DCB48F38D73F4CC6B43F34D34C",
	            INITP_02 => X"000000000000000000000000000000000000000000000000000000F00B0B0DBF",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )
	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk,
	            ADDRB => address,

DOB => instruction( 18 - 3 downto 0 ),-- OJO INSTSIZE =18
DOPB => instruction( 18 - 1 downto 18 - 2 ),-- INSTSIZE = 18
DIA => jdata( 9 - 2 downto 0 ),	 -- OJO JDATASIZE = 9
DIPA => jdata( 9 - 1 downto 9 - 1 ), -- OJO JDATASIZE = 9

	            --DOB => instruction( INSTSIZE - 3 downto 0 ),
	            --DOPB => instruction( INSTSIZE - 1 downto INSTSIZE - 2 ),
	            --DIA => jdata( JDATASIZE - 2 downto 0 ),
	            --DIPA => jdata( JDATASIZE - 1 downto JDATASIZE - 1 ),
	            
					ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	I16 : if PicoType = pbtI generate
		attribute INIT_00 of bram : label is "C00000BF00BFC00154174900501749FFC000FAA009FFF7700F20001A00EEC000" ;
		attribute INIT_01 of bram : label is "00BF00DD50234500450406004007CA01C0010AFF4017EAFF54174900501649FF" ;
		attribute INIT_02 of bram : label is "860100CE051800BA00BA00BA060100BF00BF00BF00BF00BF00BF401B860100BF" ;
		attribute INIT_03 of bram : label is "00DD052000DD052000DD052000DD05200104051000BF00BF00BF00BF542A4610" ;
		attribute INIT_04 of bram : label is "00DD052000DD052000DD053A00DD057300DD056F00DD057400DD056100DD0544" ;
		attribute INIT_05 of bram : label is "A00000DD0520A00054534610860100CE051C00BA00BA00BA00BA060100DD0520" ;
		attribute INIT_06 of bram : label is "47615874475B587347415874473A58734730157001048F010F2E5864452F15F0" ;
		attribute INIT_07 of bram : label is "408109FF5C80480AA80F187054804830A8F018700AFF00DD053F5874477B5873" ;
		attribute INIT_08 of bram : label is "090F0098408F00DD053F01048F010F2E5889452F15F0588E4C0A1C7080000900" ;
		attribute INIT_09 of bram : label is "C53040A500A6589F450A15C0010415F040811A709780070608075894270FF880" ;
		attribute INIT_0A of bram : label is "A00054ADC001000BA0000F20001A0104051000EEA0000F2F58A54F2F8F0100DD" ;
		attribute INIT_0B of bram : label is "037DA00054BBC30100B50314A00054B6C20100B00219A00054B1C10100AC0128" ;
		attribute INIT_0C of bram : label is "A4F01450A00000C4C440A4F8A000C440E40100ACC440E401A00054C0C30100B5" ;
		attribute INIT_0D of bram : label is "C40CA4F01450A000C44004F000B000CA0406040604060407145000AC00CAC408" ;
		attribute INIT_0E of bram : label is "043000BAA000C44004F000B000C4C4400406040604070407145000AC00C4C440" ;
		attribute INIT_0F of bram : label is "050100CE050C00CE050600CE052800B000CA042000B000CA00B500CA00BA00CA" ;
	begin
	    bram : component RAMB4_S8_S16
	        generic map (
	            INIT_00 => X"C00000BF00BFC00154174900501749FFC000FAA009FFF7700F20001A00EEC000",
	            INIT_01 => X"00BF00DD50234500450406004007CA01C0010AFF4017EAFF54174900501649FF",
	            INIT_02 => X"860100CE051800BA00BA00BA060100BF00BF00BF00BF00BF00BF401B860100BF",
	            INIT_03 => X"00DD052000DD052000DD052000DD05200104051000BF00BF00BF00BF542A4610",
	            INIT_04 => X"00DD052000DD052000DD053A00DD057300DD056F00DD057400DD056100DD0544",
	            INIT_05 => X"A00000DD0520A00054534610860100CE051C00BA00BA00BA00BA060100DD0520",
	            INIT_06 => X"47615874475B587347415874473A58734730157001048F010F2E5864452F15F0",
	            INIT_07 => X"408109FF5C80480AA80F187054804830A8F018700AFF00DD053F5874477B5873",
	            INIT_08 => X"090F0098408F00DD053F01048F010F2E5889452F15F0588E4C0A1C7080000900",
	            INIT_09 => X"C53040A500A6589F450A15C0010415F040811A709780070608075894270FF880",
	            INIT_0A => X"A00054ADC001000BA0000F20001A0104051000EEA0000F2F58A54F2F8F0100DD",
	            INIT_0B => X"037DA00054BBC30100B50314A00054B6C20100B00219A00054B1C10100AC0128",
	            INIT_0C => X"A4F01450A00000C4C440A4F8A000C440E40100ACC440E401A00054C0C30100B5",
	            INIT_0D => X"C40CA4F01450A000C44004F000B000CA0406040604060407145000AC00CAC408",
	            INIT_0E => X"043000BAA000C44004F000B000C4C4400406040604070407145000AC00C4C440",
	            INIT_0F => X"050100CE050C00CE050600CE052800B000CA042000B000CA00B500CA00BA00CA"
	        )
			port map (
				DIB => "0000000000000000",  
				ENB => '1', 
				WEB => '0',
				RSTB =>	'0',
				CLKB => clk,
				ADDRB => address,
				DOB => instruction( INSTSIZE - 1 downto 0 ),  
				DIA => jdata( JDATASIZE - 1 downto 0 ),   
				ENA => juser1, 
				WEA => jwrite,
				RSTA => '0',
				CLKA => clk,
				ADDRA => jaddr,
				DOA => open  
			) ; 
	end generate ;

	I20 : if PicoType = pbtS generate
		attribute INIT_00 of ram_1 : label is "3030303030333331130333033333331333310032303031313333313130000333" ;
		attribute INIT_01 of ram_1 : label is "3031003100030313131313131031031023023113033330303030303030303030" ;
		attribute INIT_02 of ram_1 : label is "0231302313023130231020330320311303331030301223100333031031031030" ;
		attribute INIT_03 of ram_1 : label is "0303030330333333032203322222033200022033222203300023202203202313" ;
		attribute INIT_04 of ram_1 : label is "0000000000000000000000000000000000000000000033000023002300312333" ;
		attribute INIT_05 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_1 : label is "3000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_2 : label is "000000000000005480000000000004800054404CC04E5454C00C5454CF0F000C" ;
		attribute INIT_01 of ram_2 : label is "4054A154A10005454545454541080541A00A5480000000000000000000000000" ;
		attribute INIT_02 of ram_2 : label is "0A5C00A5C00A5C00A5C0A00000A05480C40541014190052F0040008054154180" ;
		attribute INIT_03 of ram_2 : label is "000000000000000000AC000C0000100CCA1AC0000000100CA1A0CAACE0CEA5C0" ;
		attribute INIT_04 of ram_2 : label is "0000000000000000000000000000000000000000000045AA14A0CAA0CA52A000" ;
		attribute INIT_05 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_2 : label is "4000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_3 : label is "050505051500004660500060000000600005560A0A0A4909000049090A97F000" ;
		attribute INIT_01 of ram_3 : label is "09C8884888A0587878787878751FF85500504660500006050505050505050505" ;
		attribute INIT_02 of ram_3 : label is "304303042020410104000F01500F8FF0500855150A778878900051FF8558CC09" ;
		attribute INIT_03 of ram_3 : label is "5050505004000000400440044444400444404400444440044400440440440430" ;
		attribute INIT_04 of ram_3 : label is "0000000000000000000000000000000000000000000000878700550055150000" ;
		attribute INIT_05 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_3 : label is "1000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_4 : label is "D2D2D2D201BBBB210C1BBB0BBBBBB10BBD2000000F1F101F0BB0101F0AF721E0" ;
		attribute INIT_01 of ram_4 : label is "8F800783F7FD3777675747373700262F0D20510C1BBBB0D2D2D2D3D7D6D7D6D4" ;
		attribute INIT_02 of ram_4 : label is "70B0B10B0B10B0A20A0002101E02A20D3AA90C0F87800908098D300282F80700" ;
		attribute INIT_03 of ram_4 : label is "0C0C0C2BC2BCBCBC3B04FBC400005AC40F504FBC00005AC0F50C4F040A400C0B" ;
		attribute INIT_04 of ram_4 : label is "000000000000000000000000000000000000000000006887700CC00C80010BBC" ;
		attribute INIT_05 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_5 : label is "D0D0D0D040FFFFA01E8AAA1FFFFFFB1FFD3040711F7F706F0FF1707F00F00AE0" ;
		attribute INIT_01 of ram_5 : label is "1F0AF00000FDF4B314B314A30041E4F00D00301ECAAAA1D0D0D0DAD3DFD4D1D4" ;
		attribute INIT_02 of ram_5 : label is "D0B15406109011C80D1B00A40E0F5F1D056FA040100674F0F8FDF41E9F0EA000" ;
		attribute INIT_03 of ram_5 : label is "1ECE6E80A00A5AAA0A00004066770C40C000000A66670CA8000408001C010015" ;
		attribute INIT_04 of ram_5 : label is "00000000000000000000000000000000000000000000020F010E0F0E0FA0055E" ;
		attribute INIT_05 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_06 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_07 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_5 : label is "E000000000000000000000000000000000000000000000000000000000000000" ;

		signal data_out : std_logic_vector( 3 downto 0 ) ;
	begin
	    ram_1 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"3030303030333331130333033333331333310032303031313333313130000333",
				INIT_01 => X"3031003100030313131313131031031023023113033330303030303030303030",
				INIT_02 => X"0231302313023130231020330320311303331030301223100333031031031030",
				INIT_03 => X"0303030330333333032203322222033200022033222203300023202203202313",
				INIT_04 => X"0000000000000000000000000000000000000000000033000023002300312333",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"3000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => data_out,  
DIB => jdata( 11 downto 9 - 1 ), -- OJO JDATASIZE = 9 Y LOS DI VUELTA  ademas cambiamos el tama�o a 4 bits

				--DIB => jdata( JDATASIZE - 1 downto 16 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
			-- loose top 2 bits
			instruction( 17 downto 16 ) <= data_out( 1 downto 0 ) ;

	    ram_2 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"000000000000005480000000000004800054404CC04E5454C00C5454CF0F000C",
				INIT_01 => X"4054A154A10005454545454541080541A00A5480000000000000000000000000",
				INIT_02 => X"0A5C00A5C00A5C00A5C0A00000A05480C40541014190052F0040008054154180",
				INIT_03 => X"000000000000000000AC000C0000100CCA1AC0000000100CA1A0CAACE0CEA5C0",
				INIT_04 => X"0000000000000000000000000000000000000000000045AA14A0CAA0CA52A000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"4000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 15 downto 12 ),  
				DIB => jdata( 15 downto 12 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_3 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"050505051500004660500060000000600005560A0A0A4909000049090A97F000",
				INIT_01 => X"09C8884888A0587878787878751FF85500504660500006050505050505050505",
				INIT_02 => X"304303042020410104000F01500F8FF0500855150A778878900051FF8558CC09",
				INIT_03 => X"5050505004000000400440044444400444404400444440044400440440440430",
				INIT_04 => X"0000000000000000000000000000000000000000000000878700550055150000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"1000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 11 downto 8 ),  
				DIB => jdata( 11 downto 8 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_4 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"D2D2D2D201BBBB210C1BBB0BBBBBB10BBD2000000F1F101F0BB0101F0AF721E0",
				INIT_01 => X"8F800783F7FD3777675747373700262F0D20510C1BBBB0D2D2D2D3D7D6D7D6D4",
				INIT_02 => X"70B0B10B0B10B0A20A0002101E02A20D3AA90C0F87800908098D300282F80700",
				INIT_03 => X"0C0C0C2BC2BCBCBC3B04FBC400005AC40F504FBC00005AC0F50C4F040A400C0B",
				INIT_04 => X"000000000000000000000000000000000000000000006887700CC00C80010BBC",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 7 downto 4 ),  
				DIB => jdata( 7 downto 4 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_5 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"D0D0D0D040FFFFA01E8AAA1FFFFFFB1FFD3040711F7F706F0FF1707F00F00AE0",
				INIT_01 => X"1F0AF00000FDF4B314B314A30041E4F00D00301ECAAAA1D0D0D0DAD3DFD4D1D4",
				INIT_02 => X"D0B15406109011C80D1B00A40E0F5F1D056FA040100674F0F8FDF41E9F0EA000",
				INIT_03 => X"1ECE6E80A00A5AAA0A00004066770C40C000000A66670CA8000408001C010015",
				INIT_04 => X"00000000000000000000000000000000000000000000020F010E0F0E0FA0055E",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"E000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 3 downto 0 ),  
				DIB => jdata( 3 downto 0 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
	end generate ;

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture mix ;
